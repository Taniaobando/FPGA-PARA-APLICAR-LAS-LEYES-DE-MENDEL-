-----------------------------
--Actividad: ROM
--Autor(as): Laura Arango,Andres Salazar, Tania Obando, Verónica Tofiño.
--Fecha:15/11/2018
--Curso:Arquitectura del computador II
--
--archivo: rom.vhd
-----------------------------
--Descripcion: Memoria de dirección. Solo es de lectura
-----------------------------
--Cambios: Se añadió esta entrada.
-----------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity rom is
port (
	address: in integer range 0 to 511; -- Direcciones posibles
	data_out: out std_logic_vector (21 downto 0) -- Instrucción guardada en la ROM
);
end entity;

architecture rom_arc of rom is
signal reg_address: integer range 0 to 511; 
type memoria is array (0 to 511) of std_logic_vector(21 downto 0);
constant rom: memoria := (
0 => "0000001000000000000010", --Todas las instrucciones que usa nuestro codigo (de la 0 a la 283)
1 => "0000001100000000000001",
2 => "0000010000000000000000",
3 => "0000010100000000000011",
4 => "0000000100000000000000",
5 => "0001100100011000000000",
--5 => "0100001000001000001000",
6 => "0100001100001000001001",
7 => "0100010000001000001010",
8 => "0100010100001000001011",
9 => "1100000000000000000000",
10 => "0110001100001000000000",
11 => "1100000000000000000001",
12 => "0110010000001000000001",
13 => "1100000000000000000010",
14 => "0110010100001000000010",
15 => "1100000000000000000011",
16 => "0110011000001000000011",
17 => "1100000000000000000100",
18 => "0110011100001000000100",
19 => "1100000000000000000101",
20 => "0110100000001000000101",
21 => "1100000000000000000110",
22 => "0110100100001000000110",
23 => "1100000000000000000111",
24 => "0110101000001000000111",
25 => "0000101100000000000000",
26 => "0000110000000000000101",
27 => "0000110100000000001000",
28 => "0001011000000000000011",
29 => "0001011100000000000011",
30 => "0001100000000000000100",
31 => "0001100100000000000001",
32 => "0001101000000000000010",
33 => "0001101100000000000011",
34 => "1000101101100100011000",
35 => "0110111001101000000000",
36 => "1000111000011000101000",
37 => "0000110101101000000001",
38 => "0000101101011000000001",
39 => "1000000000000000100010",
40 => "0000110100000000001000",
41 => "0000101100000000000000",
42 => "1010101110110000101101",
43 => "1000101110111000110001",
44 => "1000101111000000101111",
45 => "0000001000000000000001",
46 => "1000000000000000110011",
47 => "0000001000000000000011",
48 => "1000000000000000110011",
49 => "0000001000000000000010",
50 => "1000000000000000110011",
51 => "1000101101100100011000",
52 => "0110111001101000000000",
53 => "1000111000111000111001",
54 => "0000110101101000000001",
55 => "0000101101011000000001",
56 => "1000000000000000110011",
57 => "0000110100000000001000",
58 => "0000101100000000000000",
59 => "1010101110110000111110",
60 => "1000101110111001000010",
61 => "1000101111000001000000",
62 => "0000111100000000000001",
63 => "1000000000000001000100",
64 => "0000111100000000000011",
65 => "1000000000000001000100",
66 => "0000111100000000000010",
67 => "1000000000000001000100",
68 => "1000101101100100011000",
69 => "0110111001101000000000",
70 => "1000111000100001001010",
71 => "0000110101101000000001",
72 => "0000101101011000000001",
73 => "1000000000000001000100",
74 => "0000110100000000001000",
75 => "0000101100000000000000",
76 => "1010101110110001001111",
77 => "1000101110111001010011",
78 => "1000101111000001010001",
79 => "0001000000000000000001",
80 => "1000000000000001010101",
81 => "0001000000000000000011",
82 => "1000000000000001010101",
83 => "0001000000000000000010",
84 => "1000000000000001010101",
85 => "1000101101100100011000",
86 => "0110111001101000000000",
87 => "1000111001000001011011",
88 => "0000110101101000000001",
89 => "0000101101011000000001",
90 => "1000000000000001010101",
91 => "0000110100000000001000",
92 => "0000101100000000000000",
93 => "1010101110110001100000",
94 => "1000101110111001100100",
95 => "1000101111000001100010",
96 => "0001000100000000000001",
97 => "1000000000000001100110",
98 => "0001000100000000000011",
99 => "1000000000000001100110",
100 => "0001000100000000000010",
101 => "1000000000000001100110",
102 => "1000101101100100011000",
103 => "0110111001101000000000",
104 => "1000111000101001101100",
105 => "0000110101101000000001",
106 => "0000101101011000000001",
107 => "1000000000000001100110",
108 => "0000110100000000001000",
109 => "0000101100000000000000",
110 => "1010101110110001110001",
111 => "1000101110111001110101",
112 => "1000101111000001110011",
113 => "0001001000000000000001",
114 => "1000000000000001110111",
115 => "0001001000000000000011",
116 => "1000000000000001110111",
117 => "0001001000000000000010",
118 => "1000000000000001110111",
119 => "1000101101100100011000",
120 => "0110111001101000000000",
121 => "1000111001001001111101",
122 => "0000110101101000000001",
123 => "0000101101011000000001",
124 => "1000000000000001110111",
125 => "0000110100000000001000",
126 => "0000101100000000000000",
127 => "1010101110110010000010",
128 => "1000101110111010000110",
129 => "1000101111000010000100",
130 => "0001001100000000000001",
131 => "1000000000000010001000",
132 => "0001001100000000000011",
133 => "1000000000000010001000",
134 => "0001001100000000000010",
135 => "1000000000000010001000",
136 => "1000101101100100011000",
137 => "0110111001101000000000",
138 => "1000111000110010001110",
139 => "0000110101101000000001",
140 => "0000101101011000000001",
141 => "1000000000000010001000",
142 => "0000110100000000001000",
143 => "0000101100000000000000",
144 => "1010101110110010010011",
145 => "1000101110111010010111",
146 => "1000101111000010010101",
147 => "0001010000000000000001",
148 => "1000000000000010011001",
149 => "0001010000000000000011",
150 => "1000000000000010011001",
151 => "0001010000000000000010",
152 => "1000000000000010011001",
153 => "1000101101100100011000",
154 => "0110111001101000000000",
155 => "1000111001010010011111",
156 => "0000110101101000000001",
157 => "0000101101011000000001",
158 => "1000000000000010011001",
159 => "0000110100000000001000",
160 => "0000101100000000000000",
161 => "1010101110110010100100",
162 => "1000101110111010101000",
163 => "1000101111000010100110",
164 => "0001010100000000000001",
165 => "0000000000000010101011",
166 => "0001010100000000000011",
167 => "0000000000000010101011",
168 => "0001010100000000000010",
169 => "0000000000000010101011",
170 => "0000110100000000000000",
171 => "1000001011001010111000",
172 => "1000001011010010111100",
173 => "1000001011011011000000",
174 => "1001000011001011000011",
175 => "1001000011010011000111",
176 => "1001000011011011001011",
177 => "1001001011001011001110",
178 => "1001001011010011010010",
179 => "1001001011011011010110",
180 => "1001010011001011011001",
181 => "1001010011010011011101",
182 => "1001010011011011100001",
183 => "1000000000000100010100",
184 => "1000111111001011100100",
185 => "1000111111010011101101",
186 => "1000111111011011100111",
187 => "1000000000000010101011",
188 => "1000111111001011101101",
189 => "1000111111010011101010",
190 => "1000111111011011100111",
191 => "1000000000000010101011",
192 => "0000001000000001100100",
193 => "0100001001101000001100",
194 => "1000000000000010101011",
195 => "1001000111001011110000",
196 => "1001000111010011111001",
197 => "1001000111011011110011",
198 => "1000000000000010101011",
199 => "1001000111001011111001",
200 => "1001000111010011110110",
201 => "1001000111011011110011",
202 => "1000000000000010101011",
203 => "0001000000000001100100",
204 => "0101000001101000001101",
205 => "1000000000000010101011",
206 => "1001001111001011111100",
207 => "1001001111010100000101",
208 => "1001001111011011111111",
209 => "1000000000000010101011",
210 => "1001001111001100000101",
211 => "1001001111010100000010",
212 => "1001001111011011111111",
213 => "1000000000000010101011",
214 => "0001001000000001100100",
215 => "0101001001101000001110",
216 => "1000000000000010101011",
217 => "1001010111001100001000",
218 => "1001010111010100010001",
219 => "1001010111011100001011",
220 => "1000000000000010101011",
221 => "1001010111001100010001",
222 => "1001010111010100001110",
223 => "1001010111011100001011",
224 => "1000000000000010101011",
225 => "0001010000000001100100",
226 => "0101010001101000001111",
227 => "1000000000000010101011",
228 => "0000001000000001001011",
229 => "0100001001101000001100",
230 => "1000000000000010101011",
231 => "0000001000000001100100",
232 => "0100001001101000001100",
233 => "1000000000000010101011",
234 => "0000001000000000000000",
235 => "0100001001101000001100",
236 => "1000000000000010101011",
237 => "0000001000000000110010",
238 => "0100110001101000001100",
239 => "1000000000000010101011",
240 => "0001000000000001001011",
241 => "0101000001101000001101",
242 => "1000000000000010101011",
243 => "0001000000000001100100",
244 => "0101000001101000001101",
245 => "1000000000000010101011",
246 => "0001000000000000000000",
247 => "0101000001101000001101",
248 => "1000000000000010101011",
249 => "0001000000000000110010",
250 => "0101000001101000001101",
251 => "1000000000000010101011",
252 => "0001001000000001001011",
253 => "0101001001101000001110",
254 => "1000000000000010101011",
255 => "0001001000000001100100",
256 => "0101001001101000001110",
257 => "1000000000000010101011",
258 => "0001001000000000000000",
259 => "0101001001101000001110",
260 => "1000000000000010101011",
261 => "0001001000000000110010",
262 => "0101001001101000001110",
263 => "1000000000000010101011",
264 => "0001010000000001001011",
265 => "0101010001101000001111",
266 => "1000000000000010101011",
267 => "0001010000000001100100",
268 => "0101010001101000001111",
269 => "1000000000000010101011",
270 => "0001010000000000000000",
271 => "0101010001101000001111",
272 => "1000000000000010101011",
273 => "0001010000000000110010",
274 => "0101010001101000001111",
275 => "1000000000000010101011",
276 => "1110000000000000001100",
277 => "1110000000000000001101",
278 => "1110000000000000001110",
279 => "1110000000000000001111",
280 => "1110000000000000001010",
281 => "1110000000000000001010",
282 => "1110000000000000001010",
283 => "1110000000000000001010",
others  => "0000000000000000000000"

);
begin
	--regristar la direción
	process (address) is
	begin
		--if MemIRead = '1' then
			reg_address <= address;
			data_out <= rom(reg_address);
		--end if;
	end process;
end architecture;